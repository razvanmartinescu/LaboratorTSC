/***********************************************************************
 * A SystemVerilog testbench for an instruction register.
 * The course labs will convert this to an object-oriented testbench
 * with constrained random test generation, functional coverage, and
 * a scoreboard for self-verification.
 **********************************************************************/

module instr_register_test  // se declara un modul(unit functionala - structura in care declaram)
  import instr_register_pkg::*;  // user-defined types are defined in instr_register_pkg.sv
  (
	tb_ifc.TB intf_lab 
  );
  
  //opcode_t -> contine semnale logice 
  //timeunit 1ns/1ns;

  int seed = 555; // val initiala de tip int, val init de unde se incepe randomizarea(se da la rand)

  initial begin //timp de simulare 0
    $display("\n\n***********************************************************"); // 
    $display(    "***  THIS IS NOT A SELF-CHECKING TESTBENCH (YET).  YOU  ***");
    $display(    "***  NEED TO VISUALLY VERIFY THAT THE OUTPUT VALUES     ***");
    $display(    "***  MATCH THE INPUT VALUES FOR EACH REGISTER LOCATION  ***");
    $display(    "***********************************************************");
    $display(    "FIRST HEADER");

    $display("\nReseting the instruction register...");
    intf_lab.cb.write_pointer  <= 5'h00;         // initialize write pointer, ia val 0 
    intf_lab.cb.read_pointer   <= 5'h1F;         // initialize read pointer, ia val 1F
    intf_lab.cb.load_en        <= 1'b0;          // initialize load control line, ia val 0 
    intf_lab.cb.reset_n       <= 1'b0;          // assert reset_n (active low), ia val 0 
    repeat (2) @(posedge intf_lab.cb.clk) ;     // asteapta 2 fronturi pozitive de ceas
    intf_lab.cb.reset_n        <= 1'b1;          // deassert reset_n (active low)

    $display("\nWriting values to register stack...");
    @(posedge intf_lab.cb.clk) intf_lab.cb.load_en <= 1'b1;  // enable writing to register
    repeat (3) begin
      @(posedge intf_lab.cb.clk) randomize_transaction; // rand_trasc = functie
      //in task se pot pune val temporare (@posde)
      //in functie nu pot pune val temp
      @(negedge intf_lab.cb.clk) print_transaction; //printeaza -> functie orint_trans
    end
    @(posedge intf_lab.cb.clk) intf_lab.cb.load_en <= 1'b0;  // turn-off writing to register

    // read back and display same three register locations
    $display("\nReading back the same register locations written...");
    for (int i=0; i<=2; i++) begin
      // later labs will replace this loop with iterating through a
      // scoreboard to determine which addresses were written and
      // the expected values to be read back
      @(posedge intf_lab.cb.clk) intf_lab.cb.read_pointer <= i;
      @(negedge intf_lab.cb.clk) print_results;
    end

    @(posedge intf_lab.cb.clk) ;
    $display("\n***********************************************************");
    $display(  "***  THIS IS NOT A SELF-CHECKING TESTBENCH (YET).  YOU  ***");
    $display(  "***  NEED TO VISUALLY VERIFY THAT THE OUTPUT VALUES     ***");
    $display(  "***  MATCH THE INPUT VALUES FOR EACH REGISTER LOCATION  ***");
    $display(  "***********************************************************\n");
    $finish;
  end

  function void randomize_transaction;
    // A later lab will replace this function with SystemVerilog
    // constrained random values
    //
    // The stactic temp variable is required in order to write to fixed
    // addresses of 0, 1 and 2.  This will be replaceed with randomizeed
    // write_pointer values in a later lab
    //
    static int temp = 0;
    intf_lab.cb.operand_a     <= $random(seed)%16;                 // between -15 and 15
    intf_lab.cb.operand_b     <= $unsigned($random)%16;            // between 0 and 15
    intf_lab.cb.opcode        <= opcode_t'($unsigned($random)%8);  // between 0 and 7, cast to opcode_t type, doar poztiv
    //opcode_t' -> operatia de cast - trece din index in string
    intf_lab.cb.write_pointer <= temp++; //temp are val 0,  
  endfunction: randomize_transaction

  function void print_transaction; //printeaza 
    $display("Writing to register location %0d: ", intf_lab.cb.write_pointer);
    $display("  opcode = %0d (%s)", intf_lab.cb.opcode, intf_lab.cb.opcode.name);
    $display("  operand_a = %0d",   intf_lab.cb.operand_a);
    $display("  operand_b = %0d", intf_lab.cb.operand_b);
    $display("PRINT TRANSACTION TIME: %t\n", $time());
  endfunction: print_transaction

  function void print_results;
    $display("Read from register location %0d: ", intf_lab.cb.read_pointer);
    $display("  opcode = %0d (%s)", intf_lab.cb.instruction_word.opc, intf_lab.cb.instruction_word.opc.name);
    $display("  operand_a = %0d",   intf_lab.cb.instruction_word.op_a);
    $display("  operand_b = %0d", intf_lab.cb.instruction_word.op_b);
    $display("PRINT TRANSACTION TIME: %t\n", $time());
  endfunction: print_results

endmodule: instr_register_test